library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity MODULE is
  port( CLK, RESET: in std_logic;
        LED0: out std_logic;
        LED1: out std_logic;
        LED2: out std_logic;
        LED3: out std_logic);
end MODULE;

architecture arch of MODULE is
--##INSERT YOUR CODE HERE 

--##INSERT YOUR CODE HERE END
end;

